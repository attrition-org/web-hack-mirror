--02:28:35--  http://www.asamblea.gob.sv:80/
           => `www.asamblea.gob.sv/index.html'
Connecting to www.asamblea.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 37 [text/html]

    0K ->                                                        [100%]

02:28:36 (36.13 KB/s) - `www.asamblea.gob.sv/index.html' saved [37/37]

Converting www.asamblea.gob.sv/index.html... done.

FINISHED --02:28:36--
Downloaded: 37 bytes in 1 files
