--02:05:32--  http://www.transexpress.com.sv:80/
           => `www.transexpress.com.sv/index.html'
Connecting to www.transexpress.com.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]

    0K ->

02:05:33 (171.88 KB/s) - `www.transexpress.com.sv/index.html' saved [176]

Converting www.transexpress.com.sv/index.html... done.

FINISHED --02:05:33--
Downloaded: 176 bytes in 1 files
