--11:21:44--  http://www.fsv.gob.sv:80/
           => `www.fsv.gob.sv/index.html'
Connecting to www.fsv.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 71 [text/html]

    0K ->                                                        [100%]

11:21:48 (1.98 KB/s) - `www.fsv.gob.sv/index.html' saved [71/71]

Converting www.fsv.gob.sv/index.html... done.

FINISHED --11:21:48--
Downloaded: 71 bytes in 1 files
