--13:31:49--  http://www.minec.gob.sv:80/
           => `www.minec.gob.sv/index.html'
Connecting to www.minec.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 184 [text/html]

    0K ->                                                        [100%]

13:31:50 (179.69 KB/s) - `www.minec.gob.sv/index.html' saved [184/184]

Converting www.minec.gob.sv/index.html... done.

FINISHED --13:31:50--
Downloaded: 184 bytes in 1 files
