--19:14:39--  http://www.ads.org.sv:80/
           => `www.ads.org.sv/index.html'
Connecting to www.ads.org.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 41 [text/html]

    0K ->                                                        [100%]

19:14:41 (40.04 KB/s) - `www.ads.org.sv/index.html' saved [41/41]

Converting www.ads.org.sv/index.html... done.

FINISHED --19:14:41--
Downloaded: 41 bytes in 1 files
