--02:17:12--  http://www.emprende.org.sv:80/
           => `www.emprende.org.sv/index.html'
Connecting to www.emprende.org.sv:80... connected!
HTTP request sent, awaiting response... 
Read error (Connection reset by peer) in headers.
Retrying.

--02:17:17--  http://www.emprende.org.sv:80/
  (try: 2) => `www.emprende.org.sv/index.html'
Connecting to www.emprende.org.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 30 [text/html]

    0K ->                                                        [100%]

02:17:19 (33.04 B/s) - `www.emprende.org.sv/index.html' saved [30/30]

Converting www.emprende.org.sv/index.html... done.

FINISHED --02:17:19--
Downloaded: 30 bytes in 1 files
