--03:01:17--  http://www.fsv.gob.sv:80/
           => `www.fsv.gob.sv/index.html'
Connecting to www.fsv.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: unspecified [text/html]

    0K ->

03:01:19 (374.02 KB/s) - `www.fsv.gob.sv/index.html' saved [383]

Converting www.fsv.gob.sv/index.html... done.

FINISHED --03:01:19--
Downloaded: 383 bytes in 1 files
Converting www.fsv.gob.sv/index.html... done.
