--13:26:41--  http://www.castaneda.com.sv:80/
           => `www.castaneda.com.sv/index.html'
Connecting to www.castaneda.com.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 778 [text/html]

    0K ->                                                        [100%]

13:26:46 (251.94 B/s) - `www.castaneda.com.sv/index.html' saved [778/778]

Converting www.castaneda.com.sv/index.html... done.

FINISHED --13:26:46--
Downloaded: 778 bytes in 1 files
