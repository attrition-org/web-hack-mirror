--11:39:19--  http://www.mccann.com.sv:80/
           => `www.mccann.com.sv/index.html'
Connecting to www.mccann.com.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 214 [text/html]

    0K ->                                                        [100%]

11:39:21 (208.98 KB/s) - `www.mccann.com.sv/index.html' saved [214/214]

Loading robots.txt; please ignore errors.
--11:39:21--  http://www.mccann.com.sv:80/no-robots.txt
           => `www.mccann.com.sv/no-robots.txt'
Connecting to www.mccann.com.sv:80... connected!
HTTP request sent, awaiting response... 404 Object Not Found
11:39:21 ERROR 404: Object Not Found.

--11:39:21--  http://www.mccann.com.sv:80/n0p1z.jpg
           => `www.mccann.com.sv/n0p1z.jpg'
Connecting to www.mccann.com.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 74,708 [image/jpeg]

    0K -> .......... .......... .......... .......... .......... [ 68%]
   50K -> .......... .......... ..                               [100%]

11:40:37 (1007.58 B/s) - `www.mccann.com.sv/n0p1z.jpg' saved [74708/74708]

Converting www.mccann.com.sv/index.html... done.

FINISHED --11:40:37--
Downloaded: 74,922 bytes in 2 files
Converting www.mccann.com.sv/index.html... done.
