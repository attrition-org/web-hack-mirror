--05:03:48--  http://www.minec.gob.sv:80/
           => `www.minec.gob.sv/index.html'
Connecting to www.minec.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 649 [text/html]

    0K ->                                                        [100%]

05:03:49 (633.79 KB/s) - `www.minec.gob.sv/index.html' saved [649/649]

Loading robots.txt; please ignore errors.
--05:03:50--  http://www.minec.gob.sv:80/no-robots.txt
           => `www.minec.gob.sv/no-robots.txt'
Connecting to www.minec.gob.sv:80... connected!
HTTP request sent, awaiting response... 404 Objeto no encontrado
05:03:51 ERROR 404: Objeto no encontrado.

--05:03:51--  http://www.minec.gob.sv:80/x-s.jpg
           => `www.minec.gob.sv/x-s.jpg'
Connecting to www.minec.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 14,897 [image/jpeg]

    0K -> .......... ....                                        [100%]

05:03:54 (8.54 KB/s) - `www.minec.gob.sv/x-s.jpg' saved [14897/14897]

--05:03:54--  http://www.minec.gob.sv:80/backup.txt
           => `www.minec.gob.sv/backup.txt'
Connecting to www.minec.gob.sv:80... connected!
HTTP request sent, awaiting response... 200 OK
Length: 12,394 [text/plain]

    0K -> .......... ..                                          [100%]

05:03:56 (9.32 KB/s) - `www.minec.gob.sv/backup.txt' saved [12394/12394]

Converting www.minec.gob.sv/index.html... done.

FINISHED --05:03:56--
Downloaded: 27,940 bytes in 3 files
Converting www.minec.gob.sv/index.html... done.
